library ieee;
use ieee.std_logic_1164.all;

Entity sll1 is
 Port (
  A : in std_logic_vector(15 downto 0);
  Y : out std_logic_vector(15 downto 0));
 End;

Architecture behavior of sll1 is
begin
 Y <= A(14 downto 0) & '0';
end;