library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_signed.all;
use ieee.numeric_std.all;
-- VHDL code for ALU of the MIPS Processor
entity ALU_VHDL is
generic(
 nr_of_bits : positive := 32
);
port(
 clk : in std_logic;
 a,b : in std_logic_vector(15 downto 0); -- src1, src2
 aluop : in std_logic_vector(2 downto 0); -- function select
 alu_result: out std_logic_vector(15 downto 0); -- ALU Output Result
 mult_high: out std_logic_vector(15 downto 0); -- multipication Output high
 mult_low: out std_logic_vector(15 downto 0); -- multipication Output low
 zero: out std_logic; -- Zero Flag
 z_flag, n_flag : out std_logic
 );
end ALU_VHDL;

architecture Behavioral of ALU_VHDL is
signal result: std_logic_vector(15 downto 0);
signal M : signed((2*nr_of_bits) downto 0) := (others => '0');
signal S : signed((2*nr_of_bits) downto 0) := (others => '0');
signal P : signed((2*nr_of_bits) downto 0) := (others => '0');
signal index : natural := 0;
begin
process(clk,aluop,a,b)
variable P_temp : signed(P'range);
begin
if rising_edge(clk) then
 case aluop is
 when "000" =>
  result <= a + b; -- add
 when "001" =>
  result <= a - b; -- sub
 when "010" => 
  result <= a and b; -- and
 when "011" =>
  result <= a or b; -- or
 when "100" =>
  result <= std_logic_vector(shift_left(unsigned(a), to_integer(unsigned(b)))); 
 when "101" => --compare
  if (a - b = 0) then
   z_flag <= '1';
  end if;
  if (a - b < 0) then
   n_flag <= '1';
  end if;
  if (a - b > 0) then
   z_flag <= '0';
   n_flag <= '0'; 
  end if;
  when "110" => --multiply
   if index = 0 then
     M((2*nr_of_bits) downto nr_of_bits+1) <= to_signed(to_integer(unsigned(a)), nr_of_bits);
     S((2*nr_of_bits) downto nr_of_bits+1) <= to_signed(-to_integer(unsigned(a)), nr_of_bits);
     P(nr_of_bits downto 1) <= to_signed(to_integer(unsigned(b)), nr_of_bits);
    elsif index < (nr_of_bits+1) then
     P_temp := P;
    if P(1 downto 0) = "01" then
     P_temp := P + M;
    elsif P(1 downto 0) = "10" then
     P_temp := P + S;
    end if;
     P <= shift_right(P_temp, 1);
   end if;
   index <= index + 1;
 when others => result <= a + b; -- add
 end case;
end if;
end process;
  zero <= '1' when result=x"0000" else '0';
  alu_result <= result;
  mult_high <= std_logic_vector(P((2*nr_of_bits) downto nr_of_bits+1));
  mult_low <= std_logic_vector(P(nr_of_bits downto 1));
end Behavioral;